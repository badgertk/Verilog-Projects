`include "config.v"
/**************************************
* Module: Fetch
* Date:2013-11-24  
* Author: isaac     
*
* Description: Master Instruction Fetch Module
***************************************/
module  IF
(
    input CLK,
    input RESET,
    //This should contain the fetched instruction
    output reg [31:0] Instr1_OUT,
    //This should contain the address of the fetched instruction [DEBUG purposes]
    output reg [31:0] Instr_PC_OUT,
    //This should contain the address of the instruction after the fetched instruction (used by ID)
    output reg [31:0] Instr_PC_Plus4,

    //Will be set to true if we need to just freeze the fetch stage.
    input STALL,
    
    //There was probably a branch -- please load the alternate PC instead of Instr_PC_Plus4.
    input Request_Alt_PC,
    //Alternate PC to load
    input [31:0] Alt_PC,
    
    //Address from which we want to fetch an instruction
     output [31:0] Instr_address_2IM,
//     //Address to use for first instruction to fetch when coming out of reset
//     input [31:0]   PC_init,
     //Instruction received from instruction memory
     input [31:0]   Instr1_fIM,
	 input delay_slot_needed,
	 input cache_miss
);

wire [31:0] IncrementAmount;


assign IncrementAmount = 32'd4; //NB: This might get modified for superscalar.
reg first_stall;
reg [31:0] delay_slot_instr;
reg [31:0] delay_slot_pc;
reg delay_slot_flag;


`ifdef INCLUDE_IF_CONTENT
assign Instr_address_2IM = (Request_Alt_PC)?Alt_PC:Instr_PC_Plus4;

`else

//assign Instr_address_2IM = Instr_PC_Plus4;  //Are you sure that this is correct?

`endif

always @(posedge CLK or negedge RESET) begin
	$display("FETCH: STALL = %x", STALL);
	$display("FETCH:Instr_address_2IM = %x?%x:%x", Request_Alt_PC, Alt_PC, Instr_PC_Plus4);
    if(delay_slot_needed && !cache_miss) begin
		delay_slot_flag <= 1;
	end
	if(!RESET) begin
        Instr1_OUT <= 0;
        Instr_PC_OUT <= 0;
        Instr_PC_Plus4 <= 32'hBFC00000;
        $display("FETCH [RESET] Fetching @%x", Instr_PC_Plus4);
    end else if(CLK) begin
        if(!STALL) begin
			if(delay_slot_flag) begin
				$display("<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<TRIGGERED>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>");
				Instr1_OUT <= delay_slot_instr;
				Instr_PC_OUT <= delay_slot_pc;
				delay_slot_flag <= 0;
			end
			else begin
						Instr1_OUT <= Instr1_fIM;
						Instr_PC_OUT <= Instr_address_2IM;
			end
			//Instr1_OUT <= Instr1_fIM;
			//Instr_PC_OUT <= Instr_address_2IM;
			first_stall <= 1;

`ifdef INCLUDE_IF_CONTENT
                Instr_PC_Plus4 <= Instr_address_2IM + IncrementAmount;
                $display("FETCH:Instr@%x=%x;Next@%x",Instr_address_2IM,Instr1_fIM,Instr_address_2IM + IncrementAmount);
`else
                /* You should probably assign something to Instr_PC_Plus4. */
				
                $display("FETCH:Instr@%x=%x;Next@%x",Instr_address_2IM,Instr1_fIM,Instr_address_2IM + IncrementAmount);
                $display("FETCH:ReqAlt[%d]=%x",Request_Alt_PC,Alt_PC);
`endif
        end else begin
            $display("FETCH: Stalling; next request will be %x",Instr_address_2IM);

			if(first_stall) begin
				$display(">>>>>>>>>>>>>>>>>>%x<<<<<<<<<<<<<<<<<<<<<<%d",Instr1_fIM,Request_Alt_PC);
				if (delay_slot_needed) begin
					delay_slot_instr <= Instr1_fIM;
					delay_slot_pc <= Instr_address_2IM;
				end
			end
			first_stall <= 0;
        end
    end
	$display("Delay Slot Needed: %d", delay_slot_needed);
	$display("FETCH: Instr1_OUT = %x @ %x", Instr1_OUT, Instr_PC_OUT);
	$display("first_stall = %b", first_stall);
	$display("delay_slot_instr = %x @ %x", delay_slot_instr, delay_slot_pc);
end

endmodule

